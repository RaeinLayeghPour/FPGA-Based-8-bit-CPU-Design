library verilog;
use verilog.vl_types.all;
entity Part2_vlg_vec_tst is
end Part2_vlg_vec_tst;
