library verilog;
use verilog.vl_types.all;
entity registerB_vlg_vec_tst is
end registerB_vlg_vec_tst;
